library verilog;
use verilog.vl_types.all;
entity attention_manager is
    generic(
        WIDTH           : integer := 8
    );
    port(
        int_a           : in     vl_logic_vector;
        s_calli         : in     vl_logic_vector;
        s_reti          : in     vl_logic_vector;
        data_a          : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of WIDTH : constant is 1;
end attention_manager;
